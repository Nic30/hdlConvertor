module top;
	clocking bus @(posedge clock1);
	default input #10ns output #2ns;
	input data, ready, enable = top.mem1.enable;
	output negedge ack;
	input #1step addr;
	endclocking
endmodule