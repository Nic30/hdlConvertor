LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
PACKAGE types IS
    TYPE TestEnum IS (TestEnum1, TestEnum2, TestEnum3);
    TYPE TestArray1DUB IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE TestArray1DUU IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR;
    TYPE TestArray1DBB IS ARRAY (7 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE TestArray1DBU IS ARRAY (7 DOWNTO 0) OF STD_LOGIC_VECTOR;
    TYPE TestArray2DUB IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE TestArray2DUU IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_LOGIC_VECTOR;
    TYPE TestArray2DBB IS ARRAY (7 DOWNTO 0, 7 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    TYPE TestArray2DBU IS ARRAY (7 DOWNTO 0, 7 DOWNTO 0) OF STD_LOGIC_VECTOR;
    TYPE TestInt IS RANGE -100 TO 100;
    TYPE TestFloat IS RANGE 1.000000e+10 TO 2.000000e+10;
    SUBTYPE TestInt2 IS TestInt RANGE 0 TO TestInt'HIGH;
    SUBTYPE TestFloat2 IS TestFloat RANGE 0.000000e+00 TO TestFloat'HIGH;
    TYPE TIME IS RANGE -2147483647 TO 2147483647
        UNITS
            fs;
            ps = 1000 fs;
            ns = 1000 ps;
            us = 1000 ns;
            ms = 1000 us;
            sec = 1000 ms;
            min = 60 sec;
            hr = 60 min;
        END UNITS;
END PACKAGE;

