class C;
rand int x;
constraint proto1;
extern constraint proto2;
endclass
