virtual class BasePacket;
pure virtual function integer send(bit[31:0] data); // No implementation
endclass
