class Demo ;
integer x;
function new (integer x);
this.x = x;
endfunction
endclass
