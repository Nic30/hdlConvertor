class Packet;
integer command;
function new();
command = IDLE;
endfunction
endclass
