package example is
 constant MAX_NLBIST 		      : natural := 128;--changed from 16;
 constant MAX_NMCUT 		      : natural := 512;--changed from 96
 constant MAX_NRAM		      : natural := 512;--changed from 96
 constant MAX_NROM		      : natural := 512;--changed from 96
 -- Defines the reset value for each register
 constant STCU_MB_CTRL_RES  : mb_res_reg 
          := (
	    X"00000000", -- Index 88
	    X"00000000", -- Index 87
            X"00000000", -- Index 86
            X"00000000", -- Index 85
            X"00000000", -- Index 84
	    X"00000000", -- Index 83
            X"00000000", -- Index 82
            X"00000000", -- Index 81
            X"00000000", -- Index 80
            X"00000000", -- Index 79
	        X"00000000", -- Index 78
            X"00000000", -- Index 77
            X"00000000", -- Index 76
            X"00000000", -- Index 75
            X"00000000", -- Index 74
	        X"00000000", -- Index 73
            X"00000000", -- Index 72
            X"00000000", -- Index 71
            X"00000000", -- Index 70
            X"00000000", -- Index 69
            X"00000000", -- Index 68
            X"00000000", -- Index 67
            X"00000000", -- Index 66
            X"00000000", -- Index 65
	        X"00000000", -- Index 64
            X"00000000", -- Index 63
            X"00000000", -- Index 62
            X"00000000", -- Index 61
	        X"00000000", -- Index 60
            X"00000000", -- Index 59
            X"00000000", -- Index 58
            X"00000000", -- Index 57
	        X"00000000", -- Index 56
            X"00000000", -- Index 55
            X"00000000", -- Index 54
            X"00000000", -- Index 53
	        X"00000000", -- Index 52
            X"00000000", -- Index 51
            X"00000000", -- Index 50
            X"00000000", -- Index 49
	        X"00000000", -- Index 48
            X"00000000", -- Index 47
            X"00000000", -- Index 46
            X"00000000", -- Index 45
            X"00000000", -- Index 44
	        X"00000000", -- Index 43
            X"00000000", -- Index 42
            X"00000000", -- Index 41
            X"00000000", -- Index 40
            X"00000000", -- Index 39
	        X"00000000", -- Index 38
            X"00000000", -- Index 37
            X"00000000", -- Index 36
            X"00000000", -- Index 35
            X"00000000", -- Index 34
            X"00000000", -- Index 33
            X"00000000", -- Index 32
            X"00000000", -- Index 31
            X"00000000", -- Index 30
	        X"00000000", -- Index 29
            X"00000000", -- Index 28
            X"00000000", -- Index 27
            X"00000000", -- Index 26
	        X"00000000", -- Index 25
            X"00000000", -- Index 24
            X"00000000", -- Index 23
            X"00000000", -- Index 22
	        X"00000000", -- Index 21
            X"00000000", -- Index 20
            X"00000000", -- Index 19
            X"00000000", -- Index 18
	        X"00000000", -- Index 17
            X"00000000", -- Index 16
            X"00000000", -- Index 15
            X"00000000", -- Index 14
	        X"00000000", -- Index 13
            X"00000000", -- Index 12
            X"00000000", -- Index 11
            X"00000000", -- Index 10
            X"00000000", -- Index 9
	        X"00000000", -- Index 8
            X"00000000", -- Index 7
            X"00000000", -- Index 6
            X"00000000", -- Index 5
            X"00000000", -- Index 4
	        X"00000000", -- Index 3
            X"00000000", -- Index 2
            X"00000000", -- Index 1
            X"00000000",	 -- Index 0
	    X"00000000", -- Index 166
            X"00000000", -- Index 165
	    X"00000000", -- Index 164
            X"00000000", -- Index 163
            X"00000000", -- Index 162
            X"00000000", -- Index 161
	    X"00000000", -- Index 160
            X"00000000", -- Index 159
            X"00000000", -- Index 158
            X"00000000", -- Index 157
	    X"00000000", -- Index 156
            X"00000000", -- Index 155
            X"00000000", -- Index 154
            X"00000000", -- Index 153
	    X"00000000", -- Index 152
            X"00000000", -- Index 151
            X"00000000", -- Index 150
            X"00000000", -- Index 149
	    X"00000000", -- Index 148
            X"00000000", -- Index 147
            X"00000000", -- Index 146
            X"00000000", -- Index 145
            X"00000000", -- Index 144
	    X"00000000", -- Index 143
            X"00000000", -- Index 142
            X"00000000", -- Index 141
            X"00000000", -- Index 140
            X"00000000", -- Index 139
            X"00000000", -- Index 138
            X"00000000", -- Index 137
            X"00000000", -- Index 136
            X"00000000", -- Index 135
	    X"00000000", -- Index 134
            X"00000000", -- Index 133
            X"00000000", -- Index 132
            X"00000000", -- Index 131
	    X"00000000", -- Index 130
            X"00000000", -- Index 129
            X"00000000", -- Index 128
            X"00000000", -- Index 127
	    X"00000000", -- Index 126
            X"00000000", -- Index 125
            X"00000000", -- Index 124
            X"00000000", -- Index 123
	    X"00000000", -- Index 122
            X"00000000", -- Index 121
            X"00000000", -- Index 120
            X"00000000", -- Index 119
	    X"00000000", -- Index 118
            X"00000000", -- Index 117
            X"00000000", -- Index 116
            X"00000000", -- Index 115
            X"00000000", -- Index 114
	    X"00000000", -- Index 113
            X"00000000", -- Index 112
            X"00000000", -- Index 111
            X"00000000", -- Index 110103+(NLBIST*NLBIST_REGS)+5+NMCUT
            X"00000000", -- Index 109
	    X"00000000", -- Index 108
            X"00000000", -- Index 107
            X"00000000", -- Index 106
            X"00000000", -- Index 105
            X"00000000", -- Index 104
            X"00000000", -- Index 103
            X"00000000", -- Index 102
            X"00000000", -- Index 101
            X"00000000", -- Index 100
	    X"00000000", -- Index 99
            X"00000000", -- Index 98
            X"00000000", -- Index 97
            X"00000000", -- Index 96
	    X"00000000", -- Index 95
            X"00000000", -- Index 94
            X"00000000", -- Index 93
            X"00000000", -- Index 92
	    X"00000000", -- Index 91
            X"00000000", -- Index 90
            X"00000000", -- Index 89
            X"00000000", -- Index 88
	    X"00000000", -- Index 87
            X"00000000", -- Index 86
            X"00000000", -- Index 85
            X"00000000", -- Index 84
	    X"00000000", -- Index 83
            X"00000000", -- Index 82
            X"00000000", -- Index 81
            X"00000000", -- Index 80
            X"00000000", -- Index 79
	        X"00000000", -- Index 78
            X"00000000", -- Index 77
            X"00000000", -- Index 76
            X"00000000", -- Index 75
            X"00000000", -- Index 74
	        X"00000000", -- Index 73
            X"00000000", -- Index 72
            X"00000000", -- Index 71
            X"00000000", -- Index 70
            X"00000000", -- Index 69
            X"00000000", -- Index 68
            X"00000000", -- Index 67
            X"00000000", -- Index 66
            X"00000000", -- Index 65
	        X"00000000", -- Index 64
            X"00000000", -- Index 63
            X"00000000", -- Index 62
            X"00000000", -- Index 61
	        X"00000000", -- Index 60
            X"00000000", -- Index 59
            X"00000000", -- Index 58
            X"00000000", -- Index 57
	        X"00000000", -- Index 56
            X"00000000", -- Index 55
            X"00000000", -- Index 54
            X"00000000", -- Index 53
	        X"00000000", -- Index 52
            X"00000000", -- Index 51
            X"00000000", -- Index 50
            X"00000000", -- Index 49
	        X"00000000", -- Index 48
            X"00000000", -- Index 47
            X"00000000", -- Index 46
            X"00000000", -- Index 45
            X"00000000", -- Index 44
	        X"00000000", -- Index 43
            X"00000000", -- Index 42
            X"00000000", -- Index 41
            X"00000000", -- Index 40
            X"00000000", -- Index 39
	        X"00000000", -- Index 38
            X"00000000", -- Index 37
            X"00000000", -- Index 36
            X"00000000", -- Index 35
            X"00000000", -- Index 34
            X"00000000", -- Index 33
            X"00000000", -- Index 32
            X"00000000", -- Index 31
            X"00000000", -- Index 30
	        X"00000000", -- Index 29
            X"00000000", -- Index 28
            X"00000000", -- Index 27
            X"00000000", -- Index 26
	        X"00000000", -- Index 25
            X"00000000", -- Index 24
            X"00000000", -- Index 23
            X"00000000", -- Index 22
	        X"00000000", -- Index 21
            X"00000000", -- Index 20
            X"00000000", -- Index 19
            X"00000000", -- Index 18
	        X"00000000", -- Index 17
            X"00000000", -- Index 16
            X"00000000", -- Index 15
            X"00000000", -- Index 14
	        X"00000000", -- Index 13
            X"00000000", -- Index 12
            X"00000000", -- Index 11
            X"00000000", -- Index 10
            X"00000000", -- Index 9
	        X"00000000", -- Index 8
            X"00000000", -- Index 7
            X"00000000", -- Index 6
            X"00000000", -- Index 5
            X"00000000", -- Index 4
	        X"00000000", -- Index 3
            X"00000000", -- Index 2
            X"00000000", -- Index 1
            X"00000000"	 -- Index 0
          );

  component demo is
    generic (
      GENERIC1: boolean := false;
      GENERIC2: integer := 100
    );
    port (
      a, b : in std_ulogic := '1';
      c, d : out std_ulogic_vector(7 downto 0);
      e, f : inout unsigned(7 downto 0)
    );
  end component;
end package;
