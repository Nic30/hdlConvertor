LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY test_entity_top IS
END ENTITY;

ARCHITECTURE test OF test_entity_top IS
    SUBTYPE DIGITS IS INTEGER RANGE 0 TO 9;
    FUNCTION RESOLVE_VALUE (SIGNAL anonymous : BIT_VECTOR) RETURN BIT;
    SUBTYPE BIT_NEW IS RESOLVE_VALUE BIT;
BEGIN
END ARCHITECTURE;
