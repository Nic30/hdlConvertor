architecture arch of module is
begin
   data <= i_data and i_mask;
end architecture arch;