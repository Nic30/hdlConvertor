architecture arch of module is
begin
    data <= i_data(i_data'range) and i_mask;
end architecture arch;