virtual class D;
pure constraint Test;
endclass
