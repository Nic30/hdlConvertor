architecture arch of module is
    signal Reg1,Reg2,Reg3 : signed(7 downto 0) := (others => '0');
begin
end architecture arch;
