`ifndef _parameters_vh_
`define _parameters_vh_
"a.vh"
`endif