module mymod (
output .P1(r[3:0]),
output .P2(r[7:4]),
ref
.Y(x),
input
R );
logic [7:0] r;
int x;
endmodule
