library IEEE;

package CONFIG is
			TYPE AddersType is (RCA, CLA, CSA, CSA_CLA);
end package ;