class vector #(parameter width = 7, type T = int);
endclass
