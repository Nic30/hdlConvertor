LIBRARY IEEE;
PACKAGE CONFIG IS
    TYPE AddersType IS (RCA, CLA, CSA, CSA_CLA);
END PACKAGE;

