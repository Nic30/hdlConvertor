covergroup zz(int bad);
cross x, y
{
illegal_bins illegal = binsof(y) intersect {bad};
}
endgroup



