class vector #(size = 1);
  logic [size-1:0] v;
endclass