package array_const_pkg is
 constant CONST_ARRAY  : externally_defined_array_t 
          := (
	    X"00000001",
	    X"00000002",
            X"00000003",
            X"00000004"
          );
end package;
