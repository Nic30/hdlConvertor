typedef int T;
class C;
extern function void f(T x);
typedef real T;
endclass
function void C::f(T x);
endfunction
