class C ;
endclass
module M #( type T = C, T p = 4,
type T2, T2 p2 = 4
) () ;
endmodule
