module top;
    real a;
    real b;
    var type((a + b)) c;
endmodule
