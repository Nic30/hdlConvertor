ARCHITECTURE arch OF module IS
BEGIN
    data <= (i_data AND i_mask);
END ARCHITECTURE;
