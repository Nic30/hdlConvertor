typedef struct {
logic [7:0] a;
bit b;
bit signed [31:0] c;
string s;
} sa;
