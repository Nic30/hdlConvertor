module top;
    real a = 4.76;
    real b = 0.74;
    var type(a + b) c;
endmodule
