`ifndef _a_vh_
`define _a_vh_
"a.vh"
`endif