ARCHITECTURE arch OF module IS
    SIGNAL Reg1 : signed(7 DOWNTO 0) := (OTHERS => '0');
    SIGNAL Reg2 : signed(7 DOWNTO 0) := (OTHERS => '0');
    SIGNAL Reg3 : signed(7 DOWNTO 0) := (OTHERS => '0');
BEGIN
END ARCHITECTURE;
