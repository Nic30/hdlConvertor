module chip;
    import chip_pkg::*;
endmodule
